netcdf tmp_jsonconvention {
dimensions:
	d1 = 1 ;
variables:
	int v(d1) ;
		v:varjson1 = "{\"key1\": [1,2,3], \"key2\": {\"key3\": \"abc\"}}" ;
		v:varjson2 = "[[1.0,0.0,0.0],[0.0,1.0,0.0],[0.0,0.0,1.0]]" ;
		v:varjson3 = "[0.,0.,1.]" ;
		v:varchar1  = "1.0, 0.0, 0.0" ;

// global attributes:
		:globalfloat = 1. ;
		:globalfloatvec = 1., 2. ;
		:globalchar = "abc" ;
		:globalillegal = "[ [ 1.0, 0.0, 0.0 ], [ 0.0, 1.0, 0.0 ], [ 0.0, 0.0, 1.0 " ;
data:

 v = _ ;
}
